library verilog;
use verilog.vl_types.all;
entity TOP_vlg_vec_tst is
end TOP_vlg_vec_tst;
